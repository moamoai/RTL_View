

module mod(
  input  [10:0] i,
  input  [12:0] i,
  output [13:0] o
);
  jkjk;
  ij
endmodule
