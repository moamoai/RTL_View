module mod(
  input  [10:0] i  [10:0],
  input  [12:0] jk [10:0][20:0],
  output [13:0] jo,
  output [13:0] o
);
  jkjk;
  ij
endmodule
